module xor8bits (S, A, B);

	output [7:0] S;
	input  [7:0] A;
	input  [7:0] B;

	// Instanciando uma porta OR para cada bit
	xor Xor0 (S[0], A[0], B[0]);
	xor Xor1 (S[1], A[1], B[1]);
	xor Xor2 (S[2], A[2], B[2]);
	xor Xor3 (S[3], A[3], B[3]);
	xor Xor4 (S[4], A[4], B[4]);
	xor Xor5 (S[5], A[5], B[5]);
	xor Xor6 (S[6], A[6], B[6]);
	xor Xor7 (S[7], A[7], B[7]);

endmodule